package regs_pkg;
  localparam logic [7:0] RegSysId0 = 8'h00;
  localparam logic [7:0] RegSysId1 = 8'h01;
  localparam logic [7:0] RegSysId2 = 8'h02;
  localparam logic [7:0] RegSysId3 = 8'h03;
  localparam logic [7:0] RegSysId4 = 8'h04;
  localparam logic [7:0] RegSysVersion = 8'h05;
endpackage


